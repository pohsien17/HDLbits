module top_module(
	input in,
	output out
);

	assign out = in ; 
	// a simple wire circuit
	
endmodule 
